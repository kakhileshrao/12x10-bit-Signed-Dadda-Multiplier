library ieee;
use ieee.std_logic_1164.all;
use work.dadda_utils.all;
use ieee.numeric_std.all;

entity dadda_multi is
  port(
    a: in std_logic_vector(9 downto 0);
    b: in std_logic_vector(11 downto 0);
    p: out std_logic_vector(21 downto 0)
  );
end dadda_multi;

architecture dadda_multi_arch of dadda_multi is
signal add_in1, add_in2 : std_logic_vector(20 downto 0);

signal l1: std_logic_vector(9 downto 0);
signal l2: std_logic_vector(9 downto 0);
signal l3: std_logic_vector(9 downto 0);
signal l4: std_logic_vector(9 downto 0);
signal l5: std_logic_vector(9 downto 0);
signal l6: std_logic_vector(9 downto 0);
signal l7: std_logic_vector(9 downto 0);
signal l8: std_logic_vector(9 downto 0);
signal l9: std_logic_vector(9 downto 0);
signal l10: std_logic_vector(9 downto 0);
signal l11: std_logic_vector(9 downto 0);
signal l12: std_logic_vector(9 downto 0);
-- Carry bits
signal c: std_logic_vector(30 downto 1);
-- Step 1
signal s1_1: std_logic_vector(20 downto 0);	
signal s1_2: std_logic_vector(18 downto 0);
signal s1_3: std_logic_vector(16 downto 0);
signal s1_4: std_logic_vector(14 downto 0);
signal s1_5: std_logic_vector(12 downto 0);
signal s1_6: std_logic_vector(10 downto 0);
signal s1_7: std_logic_vector(8 downto 0);
signal s1_8: std_logic_vector(6 downto 0);
signal s1_9: std_logic_vector(5 downto 0);
-- Step 2
signal s2_1: std_logic_vector(20 downto 0);	
signal s2_2: std_logic_vector(18 downto 0);
signal s2_3: std_logic_vector(16 downto 0);
signal s2_4: std_logic_vector(14 downto 0);
signal s2_5: std_logic_vector(12 downto 0);
signal s2_6: std_logic_vector(11 downto 0);
-- Step 3
signal s3_1: std_logic_vector(20 downto 0);	
signal s3_2: std_logic_vector(18 downto 0);
signal s3_3: std_logic_vector(16 downto 0);
signal s3_4: std_logic_vector(15 downto 0);
-- Step 4 
signal s4_1: std_logic_vector(20 downto 0);	
signal s4_2: std_logic_vector(18 downto 0);
signal s4_3: std_logic_vector(17 downto 0);
-- step 5
signal s5_1: std_logic_vector(20 downto 0);	
signal s5_2: std_logic_vector(19 downto 0);

signal C_temp,C_temp1: std_logic;


component brentkungadder_dadda is
port( a,b :in std_logic_vector(20 downto 0);
		--carry_in : in std_logic;
		--add_out: out std_logic_vector(19 downto 0));
		sum : out std_logic_vector(20 downto 0);
		carry_out : out std_logic);
		
		end component brentkungadder_dadda;

	
begin
	
	l1 <= and_8b(b(0), a); l2 <= and_8b(b(1), a);
	l3 <= and_8b(b(2), a); l4 <= and_8b(b(3), a);
	l5 <= and_8b(b(4), a); l6 <= and_8b(b(5), a);
	l7 <= and_8b(b(6), a); l8 <= and_8b(b(7), a);
	l9 <= and_8b(b(8), a); l10 <= and_8b(b(9), a);
	l11 <= and_8b(b(10), a); l12 <= and_8b2(b(11), a);


    --                      9 8  7 6 5 4 3 2 1 0
    ---------------------------------------
	-- l1                   2 * * * * * * * * *
	-- l2                 2 2 * * * * * * * * 
	-- l3               * 2 * * * * * * * *
	-- l4             * * * * * * * * * *
	-- l5           * * * * * * * * * *
	-- l6         * * * * * * * * * *
	-- l7       * * * * * * * * * *
	-- l8     * * * * * * * * * *
	-- l9   * * * * * * * * * *
    --l10 * * * * * * * * * * 

	s1_1(0) <= l1(0);
	s1_1(1) <= l1(1);
	s1_1(2) <= l1(2);
	s1_1(3) <= l1(3);
	s1_1(4) <= l1(4);
	s1_1(5) <= l1(5);
	s1_1(6) <= l1(6);
	s1_1(7) <= l1(7);
	s1_1(8) <= l1(8);
	s1_1(9) <= sum_3b(l1(9), l2(8),'1');   ---------modification done here
	s1_1(10) <= sum_3b(l2(9), l3(8), l4(7));
	s1_1(11) <= sum_3b(l3(9), l4(8), l5(7));
	s1_1(12) <= sum_3b(l4(9), l5(8), carry_2b(l12(0),'1')); --modification done here
	s1_1(13) <= l5(9);
	s1_1(14) <= l6(9);
	s1_1(15) <= l7(9);
	s1_1(16) <= l8(9);
	s1_1(17) <= l9(9);
	s1_1(18) <= l10(9);
	s1_1(19) <= l11(9);
	s1_1(20) <= l12(9);

	s1_2(0) <= l2(0);
	s1_2(1) <= l2(1);
	s1_2(2) <= l2(2);
	s1_2(3) <= l2(3);
	s1_2(4) <= l2(4);
	s1_2(5) <= l2(5);
	s1_2(6) <= l2(6);
	s1_2(7) <= l2(7);
	s1_2(8) <= l3(7);
	s1_2(9) <= l5(6);
	s1_2(10) <= l6(6);
	s1_2(11) <= l6(7);
	s1_2(12) <= l6(8);
	s1_2(13) <= l7(8);
	s1_2(14) <= l8(8);
	s1_2(15) <= l9(8);
	s1_2(16) <= l10(8);
	s1_2(17) <= l11(8);
	s1_2(18) <= l12(8);

	s1_3(0) <= l3(0);
	s1_3(1) <= l3(1);
	s1_3(2) <= l3(2);
	s1_3(3) <= l3(3);
	s1_3(4) <= l3(4);
	s1_3(5) <= l3(5);
	s1_3(6) <= l3(6);
	s1_3(7) <= l4(6);
	s1_3(8) <= l6(5);
	s1_3(9) <= l7(5);
	s1_3(10) <= l7(6);
	s1_3(11) <= l7(7);
	s1_3(12) <= l8(7);
	s1_3(13) <= l9(7);
	s1_3(14) <= l10(7);
	s1_3(15) <= l11(7);
	s1_3(16) <= l12(7);

    s1_4(0) <= l4(0);
	s1_4(1) <= l4(1);
	s1_4(2) <= l4(2);
	s1_4(3) <= l4(3);
	s1_4(4) <= l4(4);
	s1_4(5) <= l4(5);
	s1_4(6) <= l5(5);
	s1_4(7) <= l7(4);
	s1_4(8) <= l8(4);
	s1_4(9) <= l8(5);
	s1_4(10) <= l8(6);
	s1_4(11) <= l9(6);
	s1_4(12) <= l10(6);
	s1_4(13) <= l11(6);
	s1_4(14) <= l12(6);

    s1_5(0) <= l5(0);
	s1_5(1) <= l5(1);
	s1_5(2) <= l5(2);
	s1_5(3) <= l5(3);
	s1_5(4) <= l5(4);
	s1_5(5) <= l6(4);
	s1_5(6) <= l8(3);
	s1_5(7) <= l9(3);
	s1_5(8) <= l9(4);
	s1_5(9) <= l9(5);
	s1_5(10) <= l10(5);
	s1_5(11) <= l11(5);
	s1_5(12) <= l12(5);

    s1_6(0) <= l6(0);
	s1_6(1) <= l6(1);
	s1_6(2) <= l6(2);
	s1_6(3) <= l6(3);
	s1_6(4) <= l7(3);
	s1_6(5) <= l9(2);
	s1_6(6) <= l10(2);
	s1_6(7) <= l10(3);
	s1_6(8) <= l10(4);
	s1_6(9) <= l11(4);
	s1_6(10) <= l12(4);

    s1_7(0) <= l7(0);
	s1_7(1) <= l7(1);
	s1_7(2) <= l7(2);
	s1_7(3) <= l8(2);
	s1_7(4) <= l10(1);
	s1_7(5) <= l11(1);
	s1_7(6) <= l11(2);
	s1_7(7) <= l11(3);
	s1_7(8) <= l12(3);

    s1_8(0) <= l8(0);
	s1_8(1) <= l8(1);
	s1_8(2) <= l9(1);
	s1_8(3) <= l11(0);
	s1_8(4) <= sum_2b(l12(0),'1');  -- modification done here
	s1_8(5) <= l12(1);
	s1_8(6) <= l12(2);

    s1_9(0) <= l9(0);
	s1_9(1) <= l10(0);
	s1_9(2) <= carry_3b(l1(9), l2(8),'1');   ------modification done here
	s1_9(3) <= carry_3b(l2(9), l3(8), l4(7));	
	s1_9(4) <= carry_3b(l3(9), l4(8), l5(7));
	s1_9(5) <= carry_3b(l4(9), l5(8), carry_2b(l12(0),'1')); --modification done here


-- second stage-------------------------------

	s2_1(0) <= s1_1(0);
	s2_1(1) <= s1_1(1);
	s2_1(2) <= s1_1(2);
	s2_1(3) <= s1_1(3);
	s2_1(4) <= s1_1(4);
	s2_1(5) <= s1_1(5);
	s2_1(6) <= sum_2b(s1_1(6),s1_2(5));
	s2_1(7) <= sum_3b(s1_1(7),s1_2(6),s1_3(5));
	s2_1(8) <= sum_3b(s1_1(8),s1_2(7),s1_3(6));
	s2_1(9) <= sum_3b(s1_1(9),s1_2(8),s1_3(7));
	s2_1(10) <= sum_3b(s1_1(10),s1_2(9),s1_3(8));
	s2_1(11) <= sum_3b(s1_1(11),s1_2(10),s1_3(9));
	s2_1(12) <= sum_3b(s1_1(12),s1_2(11),s1_3(10));
	s2_1(13) <= sum_3b(s1_1(13),s1_2(12),s1_3(11));
	s2_1(14) <= sum_3b(s1_1(14),s1_2(13),s1_3(12));
	s2_1(15) <= sum_3b(s1_1(15),s1_2(14),s1_3(13));
	s2_1(16) <= s1_1(16);
	s2_1(17) <= s1_1(17);
	s2_1(18) <= s1_1(18);
	s2_1(19) <= s1_1(19);
	s2_1(20) <= s1_1(20);

	s2_2(0) <= s1_2(0);
	s2_2(1) <= s1_2(1);
	s2_2(2) <= s1_2(2);
	s2_2(3) <= s1_2(3);
	s2_2(4) <= s1_2(4);
	s2_2(5) <= s1_3(4);
	s2_2(6) <= sum_2b(s1_4(4),s1_5(3));
	s2_2(7) <= sum_3b(s1_4(5),s1_5(4),s1_6(3));
	s2_2(8) <= sum_3b(s1_4(6),s1_5(5),s1_6(4));
	s2_2(9) <= sum_3b(s1_4(7),s1_5(6),s1_6(5));
	s2_2(10) <= sum_3b(s1_4(8),s1_5(7),s1_6(6));
	s2_2(11) <= sum_3b(s1_4(9),s1_5(8),s1_6(7));
	s2_2(12) <= sum_3b(s1_4(10),s1_5(9),s1_6(8));
	s2_2(13) <= sum_3b(s1_4(11),s1_5(10),s1_6(9));
	s2_2(14) <= s1_4(12);
	s2_2(15) <= s1_2(15);
	s2_2(16) <= s1_2(16);
	s2_2(17) <= s1_2(17);
	s2_2(18) <= s1_2(18);

	s2_3(0) <= s1_3(0);
	s2_3(1) <= s1_3(1);
	s2_3(2) <= s1_3(2);
	s2_3(3) <= s1_3(3);
	s2_3(4) <= s1_4(3);
	s2_3(5) <= s1_6(2);
	s2_3(6) <= sum_2b(s1_7(2),s1_8(1));
	s2_3(7) <= sum_3b(s1_7(3),s1_8(2),s1_9(1));
	s2_3(8) <= sum_3b(s1_7(4),s1_8(3),s1_9(2));
	s2_3(9) <= sum_3b(s1_7(5),s1_8(4),s1_9(3));
    s2_3(10) <= sum_3b(s1_7(6),s1_8(5),s1_9(4));
    s2_3(11) <= sum_3b(s1_7(7),s1_8(6),s1_9(5));
	s2_3(12) <= s1_7(8);
	s2_3(13) <= s1_5(11);
	s2_3(14) <= s1_3(14);
	s2_3(15) <= s1_3(15);
	s2_3(16) <= s1_3(16);

	s2_4(0) <= s1_4(0);
	s2_4(1) <= s1_4(1);
	s2_4(2) <= s1_4(2);
	s2_4(3) <= s1_5(2);
	s2_4(4) <= s1_7(1);
	s2_4(5) <= s1_9(0);
	s2_4(6) <= carry_3b(s1_1(8),s1_2(7),s1_3(6));
	s2_4(7) <= carry_3b(s1_1(9),s1_2(8),s1_3(7));
	s2_4(8) <= carry_3b(s1_1(10),s1_2(9),s1_3(8));
	s2_4(9) <= carry_3b(s1_1(11),s1_2(10),s1_3(9));
	s2_4(10) <= carry_3b(s1_1(12),s1_2(11),s1_3(10));
    s2_4(11) <= carry_3b(s1_1(13),s1_2(12),s1_3(11));
	s2_4(12) <= s1_6(10);
	s2_4(13) <= s1_4(13);
	s2_4(14) <= s1_4(14);

	s2_5(0) <= s1_5(0);
	s2_5(1) <= s1_5(1);
	s2_5(2) <= s1_6(1);
	s2_5(3) <= s1_8(0);
	s2_5(4) <= carry_3b(s1_1(7),s1_2(6),s1_3(5));
	s2_5(5) <= carry_3b(s1_4(5),s1_5(4),s1_6(3));
	s2_5(6) <= carry_3b(s1_4(6),s1_5(5),s1_6(4));
	s2_5(7) <= carry_3b(s1_4(7),s1_5(6),s1_6(5));
	s2_5(8) <= carry_3b(s1_4(8),s1_5(7),s1_6(6));
	s2_5(9) <= carry_3b(s1_4(9),s1_5(8),s1_6(7)); ----------------------------------------
    s2_5(10) <= carry_3b(s1_4(10),s1_5(9),s1_6(8));
    s2_5(11) <= carry_3b(s1_1(14),s1_2(13),s1_3(12));
	s2_5(12) <= s1_5(12);

	s2_6(0) <= s1_6(0);
	s2_6(1) <= s1_7(0);
	s2_6(2) <= carry_2b(s1_1(6),s1_2(5)); --c1
	s2_6(3) <= carry_2b(s1_4(4),s1_5(3)); --c3
	s2_6(4) <= carry_2b(s1_7(2),s1_8(1)); --c6
	s2_6(5) <= carry_3b(s1_7(3),s1_8(2),s1_9(1)); --c9
	s2_6(6) <= carry_3b(s1_7(4),s1_8(3),s1_9(2)); --c12
	s2_6(7) <= carry_3b(s1_7(5),s1_8(4),s1_9(3)); --c15
	s2_6(8) <= carry_3b(s1_7(6),s1_8(5),s1_9(4)); --c18
	s2_6(9) <= carry_3b(s1_7(7),s1_8(6),s1_9(5)); --c21
	s2_6(10) <= carry_3b(s1_4(11),s1_5(10),s1_6(9)); --c23
	s2_6(11) <= carry_3b(s1_1(15),s1_2(14),s1_3(13)); --c24


-- third stage-------------------------------	

	s3_1(0) <= s2_1(0);
	s3_1(1) <= s2_1(1);
	s3_1(2) <= s2_1(2);
	s3_1(3) <= s2_1(3);
	s3_1(4) <= sum_2b(s2_1(4),s2_2(3)); --s1
	s3_1(5) <= sum_3b(s2_1(5),s2_2(4),s2_3(3)); --s2
	s3_1(6) <= sum_3b(s2_1(6),s2_2(5),s2_3(4)); --s4
	s3_1(7) <= sum_3b(s2_1(7),s2_2(6),s2_3(5)); --s6
	s3_1(8) <= sum_3b(s2_1(8),s2_2(7),s2_3(6)); --s8
	s3_1(9) <= sum_3b(s2_1(9),s2_2(8),s2_3(7)); --s10
	s3_1(10) <= sum_3b(s2_1(10),s2_2(9),s2_3(8)); --s12
	s3_1(11) <= sum_3b(s2_1(11),s2_2(10),s2_3(9)); --s14
	s3_1(12) <= sum_3b(s2_1(12),s2_2(11),s2_3(10)); --s16
	s3_1(13) <= sum_3b(s2_1(13),s2_2(12),s2_3(11)); --s18
	s3_1(14) <= sum_3b(s2_1(14),s2_2(13),s2_3(12)); --s20
	s3_1(15) <= sum_3b(s2_1(15),s2_2(14),s2_3(13)); --s22
	s3_1(16) <= sum_3b(s2_1(16),s2_2(15),s2_3(14)); --s23
    s3_1(17) <= sum_3b(s2_1(17),s2_2(16),s2_3(15)); --s24
	s3_1(18) <= s2_1(18);
	s3_1(19) <= s2_1(19);
	s3_1(20) <= s2_1(20);

	s3_2(0) <= s2_2(0);
	s3_2(1) <= s2_2(1);
	s3_2(2) <= s2_2(2);
	s3_2(3) <= s2_3(2);
	s3_2(4) <= sum_2b(s2_4(2),s2_5(1)); --s3
	s3_2(5) <= sum_3b(s2_4(3),s2_5(2),s2_6(1)); --s5
	s3_2(6) <= sum_3b(s2_4(4),s2_5(3),s2_6(2)); --s7
	s3_2(7) <= sum_3b(s2_4(5),s2_5(4),s2_6(3)); --s9
	s3_2(8) <= sum_3b(s2_4(6),s2_5(5),s2_6(4)); --s11
	s3_2(9) <= sum_3b(s2_4(7),s2_5(6),s2_6(5)); --s13
	s3_2(10) <= sum_3b(s2_4(8),s2_5(7),s2_6(6)); --s15
	s3_2(11) <= sum_3b(s2_4(9),s2_5(8),s2_6(7)); --s17
	s3_2(12) <= sum_3b(s2_4(10),s2_5(9),s2_6(8)); --s19
	s3_2(13) <= sum_3b(s2_4(11),s2_5(10),s2_6(9)); --s21
    s3_2(14) <= sum_3b(s2_4(12),s2_5(11),s2_6(10)); --s22
    s3_2(15) <= sum_3b(s2_4(13),s2_5(12),s2_6(11)); --s22
	s3_2(16) <= s2_4(14);
	s3_2(17) <= s2_2(17);
	s3_2(18) <= s2_2(18);

	s3_3(0) <= s2_3(0);
	s3_3(1) <= s2_3(1);
	s3_3(2) <= s2_4(1);
	s3_3(3) <= s2_6(0);
	s3_3(4) <= carry_3b(s2_1(5),s2_2(4),s2_3(3)); --c2
	s3_3(5) <= carry_3b(s2_1(6),s2_2(5),s2_3(4)); --c4
	s3_3(6) <= carry_3b(s2_1(7),s2_2(6),s2_3(5)); --c6
	s3_3(7) <= carry_3b(s2_1(8),s2_2(7),s2_3(6)); --c8
	s3_3(8) <= carry_3b(s2_1(9),s2_2(8),s2_3(7)); --c10
	s3_3(9) <= carry_3b(s2_1(10),s2_2(9),s2_3(8)); --c12
	s3_3(10) <= carry_3b(s2_1(11),s2_2(10),s2_3(9)); --c14
	s3_3(11) <= carry_3b(s2_1(12),s2_2(11),s2_3(10)); --c16
	s3_3(12) <= carry_3b(s2_1(13),s2_2(12),s2_3(11)); --c18
	s3_3(13) <= carry_3b(s2_1(14),s2_2(13),s2_3(12)); --c20
    s3_3(14) <= carry_3b(s2_1(15),s2_2(14),s2_3(13)); --c21
    s3_3(15) <= carry_3b(s2_1(16),s2_2(15),s2_3(14)); --c21
	s3_3(16) <= s2_3(16);

	s3_4(0) <= s2_4(0);
	s3_4(1) <= s2_5(0);
	s3_4(2) <= carry_2b(s2_1(4),s2_2(3));
	s3_4(3) <= carry_2b(s2_4(2),s2_5(1));
	s3_4(4) <= carry_3b(s2_4(3),s2_5(2),s2_6(1));
	s3_4(5) <= carry_3b(s2_4(4),s2_5(3),s2_6(2));
	s3_4(6) <= carry_3b(s2_4(5),s2_5(4),s2_6(3));
	s3_4(7) <= carry_3b(s2_4(6),s2_5(5),s2_6(4));
	s3_4(8) <= carry_3b(s2_4(7),s2_5(6),s2_6(5));
	s3_4(9) <= carry_3b(s2_4(8),s2_5(7),s2_6(6));
	s3_4(10) <= carry_3b(s2_4(9),s2_5(8),s2_6(7));
	s3_4(11) <= carry_3b(s2_4(10),s2_5(9),s2_6(8));
	s3_4(12) <= carry_3b(s2_4(11),s2_5(10),s2_6(9));
    s3_4(13) <= carry_3b(s2_4(12),s2_5(11),s2_6(10));
    s3_4(14) <= carry_3b(s2_4(13),s2_5(12),s2_6(11));
	s3_4(15) <= carry_3b(s2_1(17),s2_2(16),s2_3(15));


	-- fourth stage-------------------------------

	s4_1(0) <= s3_1(0);
	s4_1(1) <= s3_1(1);
	s4_1(2) <= s3_1(2);
	s4_1(3) <= sum_2b(s3_1(3),s3_2(2));
	s4_1(4) <= sum_3b(s3_1(4),s3_2(3),s3_3(2));
	s4_1(5) <= sum_3b(s3_1(5),s3_2(4),s3_3(3));
	s4_1(6) <= sum_3b(s3_1(6),s3_2(5),s3_3(4));
	s4_1(7) <= sum_3b(s3_1(7),s3_2(6),s3_3(5));
 	s4_1(8) <= sum_3b(s3_1(8),s3_2(7),s3_3(6));
	s4_1(9) <= sum_3b(s3_1(9),s3_2(8),s3_3(7));
	s4_1(10) <= sum_3b(s3_1(10),s3_2(9),s3_3(8));
	s4_1(11) <= sum_3b(s3_1(11),s3_2(10),s3_3(9));
	s4_1(12) <= sum_3b(s3_1(12),s3_2(11),s3_3(10));
	s4_1(13) <= sum_3b(s3_1(13),s3_2(12),s3_3(11));
	s4_1(14) <= sum_3b(s3_1(14),s3_2(13),s3_3(12));
	s4_1(15) <= sum_3b(s3_1(15),s3_2(14),s3_3(13));
	s4_1(16) <= sum_3b(s3_1(16),s3_2(15),s3_3(14));
    s4_1(17) <= sum_3b(s3_1(17),s3_2(16),s3_3(15));
    s4_1(18) <= sum_3b(s3_1(18),s3_2(17),s3_3(16));
	s4_1(19) <= s3_1(19);
	s4_1(20) <= s3_1(20);

	s4_2(0) <= s3_2(0);
	s4_2(1) <= s3_2(1);
	s4_2(2) <= s3_3(1);
	s4_2(3) <= s3_4(1);
	s4_2(4) <= s3_4(2);
	s4_2(5) <= s3_4(3);
	s4_2(6) <= s3_4(4);
	s4_2(7) <= s3_4(5);
 	s4_2(8) <= s3_4(6);
	s4_2(9) <= s3_4(7);
	s4_2(10) <= s3_4(8);
	s4_2(11) <= s3_4(9);
	s4_2(12) <= s3_4(10);
	s4_2(13) <= s3_4(11);
	s4_2(14) <= s3_4(12);
	s4_2(15) <= s3_4(13);
    s4_2(16) <= s3_4(14);
    s4_2(17) <= s3_4(15);
	s4_2(18) <= s3_2(18);

	s4_3(0) <= s3_3(0);
	s4_3(1) <= S3_4(0);
	s4_3(2) <= carry_2b(s3_1(3),s3_2(2));
	s4_3(3) <= carry_3b(s3_1(4),s3_2(3),s3_3(2));
	s4_3(4) <= carry_3b(s3_1(5),s3_2(4),s3_3(3));
	s4_3(5) <= carry_3b(s3_1(6),s3_2(5),s3_3(4));
	s4_3(6) <= carry_3b(s3_1(7),s3_2(6),s3_3(5));
	s4_3(7) <= carry_3b(s3_1(8),s3_2(7),s3_3(6));
	s4_3(8) <= carry_3b(s3_1(9),s3_2(8),s3_3(7));
	s4_3(9) <= carry_3b(s3_1(10),s3_2(9),s3_3(8));
	s4_3(10) <= carry_3b(s3_1(11),s3_2(10),s3_3(9));
	s4_3(11) <= carry_3b(s3_1(12),s3_2(11),s3_3(10));
	s4_3(12) <= carry_3b(s3_1(13),s3_2(12),s3_3(11));
	s4_3(13) <= carry_3b(s3_1(14),s3_2(13),s3_3(12));
	s4_3(14) <= carry_3b(s3_1(15),s3_2(14),s3_3(13));
	s4_3(15) <= carry_3b(s3_1(16),s3_2(15),s3_3(14));
	s4_3(16) <= carry_3b(s3_1(17),s3_2(16),s3_3(15));
	s4_3(17) <= carry_3b(s3_1(18),s3_2(17),s3_3(16));


	-- fifth stage-------------------------------

	s5_1(0) <= s4_1(0);
	s5_1(1) <= s4_1(1);
	s5_1(2) <= sum_2b(s4_1(2),s4_2(1));
	s5_1(3) <= sum_3b(s4_1(3),s4_2(2),s4_3(1)); 
	s5_1(4) <= sum_3b(s4_1(4),s4_2(3),s4_3(2)); 
	s5_1(5) <= sum_3b(s4_1(5),s4_2(4),s4_3(3)); 
	s5_1(6) <= sum_3b(s4_1(6),s4_2(5),s4_3(4)); 
	s5_1(7) <= sum_3b(s4_1(7),s4_2(6),s4_3(5)); 
	s5_1(8) <= sum_3b(s4_1(8),s4_2(7),s4_3(6)); 
	s5_1(9) <= sum_3b(s4_1(9),s4_2(8),s4_3(7)); 
	s5_1(10) <= sum_3b(s4_1(10),s4_2(9),s4_3(8)); 
	s5_1(11) <= sum_3b(s4_1(11),s4_2(10),s4_3(9)); 
	s5_1(12) <= sum_3b(s4_1(12),s4_2(11),s4_3(10)); 
	s5_1(13) <= sum_3b(s4_1(13),s4_2(12),s4_3(11)); 
	s5_1(14) <= sum_3b(s4_1(14),s4_2(13),s4_3(12)); 
	s5_1(15) <= sum_3b(s4_1(15),s4_2(14),s4_3(13)); 
	s5_1(16) <= sum_3b(s4_1(16),s4_2(15),s4_3(14)); 
	s5_1(17) <= sum_3b(s4_1(17),s4_2(16),s4_3(15)); 
	s5_1(18) <= sum_3b(s4_1(18),s4_2(17),s4_3(16)); 
    s5_1(19) <= sum_3b(s4_1(19),s4_2(18),s4_3(17)); 
	s5_1(20) <= s4_1(20); 

	s5_2(0) <= s4_2(0);
	s5_2(1) <= s4_3(0);
	s5_2(2) <= carry_2b(s4_1(2),s4_2(1));
	s5_2(3) <= carry_3b(s4_1(3),s4_2(2),s4_3(1)); 
	s5_2(4) <= carry_3b(s4_1(4),s4_2(3),s4_3(2)); 
	s5_2(5) <= carry_3b(s4_1(5),s4_2(4),s4_3(3)); 
	s5_2(6) <= carry_3b(s4_1(6),s4_2(5),s4_3(4)); 
	s5_2(7) <= carry_3b(s4_1(7),s4_2(6),s4_3(5)); 
	s5_2(8) <= carry_3b(s4_1(8),s4_2(7),s4_3(6)); 
	s5_2(9) <= carry_3b(s4_1(9),s4_2(8),s4_3(7)); 
	s5_2(10) <= carry_3b(s4_1(10),s4_2(9),s4_3(8)); 
	s5_2(11) <= carry_3b(s4_1(11),s4_2(10),s4_3(9)); 
	s5_2(12) <= carry_3b(s4_1(12),s4_2(11),s4_3(10)); 
	s5_2(13) <= carry_3b(s4_1(13),s4_2(12),s4_3(11)); 
	s5_2(14) <= carry_3b(s4_1(14),s4_2(13),s4_3(12)); 
	s5_2(15) <= carry_3b(s4_1(15),s4_2(14),s4_3(13)); 
	s5_2(16) <= carry_3b(s4_1(16),s4_2(15),s4_3(14)); 
	s5_2(17) <= carry_3b(s4_1(17),s4_2(16),s4_3(15));
	s5_2(18) <= carry_3b(s4_1(18),s4_2(17),s4_3(16));  
	s5_2(19) <= carry_3b(s4_1(19),s4_2(18),s4_3(17));

	p(0) <= s5_1(0);
	add_in1 <= '1' & s5_1(20 downto 1);
	add_in2 <= '0' & s5_2;
	Fin_add: brentkungadder_dadda port map (add_in1, add_in2, p(21 downto 1), C_temp);

end architecture;